module cache(input clk
    input [15:1] raddr0_, output reg [15:0] rdata0_, output rvalid0_,
    input [15:1] raddr1_, output reg [15:0] rdata1_, output rvalid1_,
    input wen0, input [15:1] waddr0, input [15:0] wdata0);

    parameter DELAY = 1;

    


endmodule