
module load_store_unit(
    input clk, input flush,
    
);


endmodule